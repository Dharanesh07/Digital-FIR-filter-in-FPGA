module transposed_fir #(
    parameter DATA_WIDTH = 16,
    parameter TAP_WIDTH  = 16,
    parameter TAP_COUNT  = 8
) (
    input wire i_clk,
    input wire i_rstn,
    input wire signed [DATA_WIDTH-1:0] i_fir_datain,
    output reg signed [(2*DATA_WIDTH)-1:0] o_fir_dataout,
    output reg o_fifo_wren,
    input wire sig_comp
);


  parameter ACC_WIDTH = 2 * DATA_WIDTH;

  // Coefficients and delay registers
  reg signed [TAP_WIDTH-1:0] coeff[TAP_COUNT-1:0];
  integer i, k;
  reg wren_pipeline = 1'b0;
  reg signed [(ACC_WIDTH-1):0] data_pipeline;
  reg signed [(ACC_WIDTH-1):0] acc[TAP_COUNT-1:0];
  // Load coefficients from file (if needed)



  initial begin
    for (i = 0; i < TAP_COUNT; i = i + 1) begin
      acc[i] = 0;
    end
  end

  // Transposed FIR logic
  always @(posedge i_clk) begin
    if (!i_rstn) begin
      // Reset accumulators
      coeff[0]  <= 32'b00000000000001010111000010000010;
      coeff[1]  <= 32'b00000000000001111111101010100000;
      coeff[2]  <= 32'b00000000000010100101011010011011;
      coeff[3]  <= 32'b00000000000011000000001001101101;
      coeff[4]  <= 32'b00000000000011000110011100010111;
      coeff[5]  <= 32'b00000000000010101110100101101000;
      coeff[6]  <= 32'b00000000000001101111001001100011;
      coeff[7]  <= 32'b00000000000000000000000000000000;
      coeff[8]  <= 32'b11111111111101011011101000101100;
      coeff[9]  <= 32'b11111111111010000000101111101101;
      coeff[10] <= 32'b11111111110101110001111100110110;
      coeff[11] <= 32'b11111111110000111000011011010011;
      coeff[12] <= 32'b11111111101011100001110011011110;
      coeff[13] <= 32'b11111111100110000001101111101011;
      coeff[14] <= 32'b11111111100000110000000110101000;
      coeff[15] <= 32'b11111111011100000111111000010111;
      coeff[16] <= 32'b11111111011000100100110111010011;
      coeff[17] <= 32'b11111111010110100011000110100101;
      coeff[18] <= 32'b11111111010110011010011100111011;
      coeff[19] <= 32'b11111111011000011101010000110000;
      coeff[20] <= 32'b11111111011100110111010101000011;
      coeff[21] <= 32'b11111111100011101010011111001110;
      coeff[22] <= 32'b11111111101100101110010110011011;
      coeff[23] <= 32'b11111111110111110000100100001111;
      coeff[24] <= 32'b00000000000100010100110100101111;
      coeff[25] <= 32'b00000000010001110110101011111001;
      coeff[26] <= 32'b00000000011111101010010111111000;
      coeff[27] <= 32'b00000000101101000010000000101110;
      coeff[28] <= 32'b00000000111001001101101000001010;
      coeff[29] <= 32'b00000001000011100001011100011010;
      coeff[30] <= 32'b00000001001011010110111011001110;
      coeff[31] <= 32'b00000001010000010000001100000000;
      coeff[32] <= 32'b00000001010001111010111000010100;
      coeff[33] <= 32'b00000001010000010000001100000000;
      coeff[34] <= 32'b00000001001011010110111011001110;
      coeff[35] <= 32'b00000001000011100001011100011010;
      coeff[36] <= 32'b00000000111001001101101000001010;
      coeff[37] <= 32'b00000000101101000010000000101110;
      coeff[38] <= 32'b00000000011111101010010111111000;
      coeff[39] <= 32'b00000000010001110110101011111001;
      coeff[40] <= 32'b00000000000100010100110100101111;
      coeff[41] <= 32'b11111111110111110000100100001111;
      coeff[42] <= 32'b11111111101100101110010110011011;
      coeff[43] <= 32'b11111111100011101010011111001110;
      coeff[44] <= 32'b11111111011100110111010101000011;
      coeff[45] <= 32'b11111111011000011101010000110000;
      coeff[46] <= 32'b11111111010110011010011100111011;
      coeff[47] <= 32'b11111111010110100011000110100101;
      coeff[48] <= 32'b11111111011000100100110111010011;
      coeff[49] <= 32'b11111111011100000111111000010111;
      coeff[50] <= 32'b11111111100000110000000110101000;
      coeff[51] <= 32'b11111111100110000001101111101011;
      coeff[52] <= 32'b11111111101011100001110011011110;
      coeff[53] <= 32'b11111111110000111000011011010011;
      coeff[54] <= 32'b11111111110101110001111100110110;
      coeff[55] <= 32'b11111111111010000000101111101101;
      coeff[56] <= 32'b11111111111101011011101000101100;
      coeff[57] <= 32'b00000000000000000000000000000000;
      coeff[58] <= 32'b00000000000001101111001001100011;
      coeff[59] <= 32'b00000000000010101110100101101000;
      coeff[60] <= 32'b00000000000011000110011100010111;
      coeff[61] <= 32'b00000000000011000000001001101101;
      coeff[62] <= 32'b00000000000010100101011010011011;
      coeff[63] <= 32'b00000000000001111111101010100000;
      coeff[64] <= 32'b00000000000001010111000010000010;


      for (i = 0; i < TAP_COUNT; i = i + 1) begin
        acc[i] <= 0;
      end
      o_fifo_wren   <= 1'b0;
      o_fir_dataout <= 0;
      data_pipeline <= 0;
    end else begin
      // Broadcast input to all multipliers and accumulate
        acc[0] <= i_fir_datain * coeff[0];
        for (k = 1; k < TAP_COUNT; k = k + 1) begin
          acc[k] <= acc[k-1] + (i_fir_datain * coeff[k]);
        end
        // Output the final accumulated value
        data_pipeline <= acc[TAP_COUNT-1];
        //data_pipeline <= i_fir_datain;
        // stall one clock cycle
        wren_pipeline <= 1'b1;

        o_fifo_wren   <= (wren_pipeline & (~sig_comp));
        o_fir_dataout <= data_pipeline;
    end
  end

endmodule

